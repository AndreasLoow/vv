module final_nonblocking;

logic a;

// Has no effect
final a <= 0;

endmodule
