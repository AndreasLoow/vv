module display_empty2;

initial $display("foo",,"bar");

endmodule
