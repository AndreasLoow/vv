module var_net;

logic a;

wire a;
   
endmodule
