module final_delay;

logic a;

final #1 a = 1;

endmodule
