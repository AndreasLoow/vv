module finish_finish;

initial $finish(0);

final $finish(1);

endmodule
