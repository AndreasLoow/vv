module net_init4;

wire a;

// Suspicious cycle, results in "a" being x in
// simulators, which could be a little surprising

assign a = a;

initial $monitor("a = %b for time %d", a, $time);

endmodule
