module empty_delay1;

// Edge-case

initial #1;
   
always #1;

endmodule
