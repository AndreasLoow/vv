// Unnamed example, p. 91--92

module ex4_nondet;

// MOD: rega not declared in original example since
//      just code snippet
logic rega;

initial #5 rega = 1'b1;

initial #5 rega = 1'b0;

initial #6 $display("rega at time = %d is %b", $time, rega);

/* The above may result in 1 or 0 depending on the simulation run and the simulator tool */

endmodule
