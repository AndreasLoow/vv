module cont_var4;

logic a;

assign a = 0;

assign a = 1;

endmodule
