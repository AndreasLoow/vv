module readme;

// The modules in this directory discusses
// Chen et al.'s OOPSLA'23 paper
// "The Essence of Verilog: A Tractable and Tested
// Operational Semantics for Verilog".

// The ex521 modules are inspired by the 
// example "5.1.2 Hidden Data-races"
// and private communication with the authors.

endmodule
