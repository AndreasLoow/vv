module empty;

// See the modules under 00 in the top-left menu for
// some introductory notes on how to use VV and
// notes on the semantics of Verilog.

// The other modules included illustrate various
// aspects of the semantics Verilog. The modules are
// commented and grouped by theme, e.g., modules
// discussing continuous assignments can be found
// under "cont" and modules discussing final blocks
// can be found under "end".

// See https://github.com/AndreasLoow/vv for more
// information.

endmodule
