module final2;

logic a;

initial $finish;

final a = 0;

endmodule
