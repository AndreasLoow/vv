module always_comb_writes_removed;

// variables written to be always_comb are removed
// from sensitivity list

logic a, b, c, d;

// does not include a
always_comb begin
 a = 0;
 b = a;
end

// does not include c
always_comb begin
 d = c;
 c = 0;
end

endmodule
