module net_init2;

// Page 98 of the standard says:
// "The default initialization value for a net
// shall be the value z."
//
// Based on the above the above one might maybe
// expect that the below should be able to print
// z or 0.

wire a;

assign a = 0;

initial $display("%b", a);

// However, some simulators print x here.
//
// One way to make sense of this is that the
// resolution function of the net is run before
// the drivers are initialised.

// In VV, we simply assign z as the initial value
// for unconnected nets and x as the initial value
// for connected nets, modelling a run of the
// resolution function of the net at initialisation.

endmodule
