module readme;

// The modules in this directory are based on the some of the
// issues with the Verilog standard raised in
// Documentation/developer/guide/misc/ieee1364-notes.rst
// from the Icarus Verilog simulator: https://github.com/steve/iverilog.
//
// The modules here are based on ieee1364-notes.rst from Git commit 9e4c4d5
//
// Note that ieee1364-notes.rst discusses legacy versions of the Verilog
// standard, not the latest version.

endmodule
