module wait1;

logic v;
   
initial wait(v) v = 0;

initial v = 1;

endmodule
