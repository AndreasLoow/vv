module always_comb_delay2;

logic a;

always_comb a = #1 1;

endmodule
