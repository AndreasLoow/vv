module var_var;

logic a;

logic a;

endmodule
