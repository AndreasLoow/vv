module cont_var2;

logic a;

always @(*) a = 0;

// Mixed types of assignments not allowed
assign a = 1;

endmodule
