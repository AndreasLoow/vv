module var_init1;

// Initialisation of variables is a little trick in
// Verilog because of the history of the language.
// That is, different versions of Verilog handle
// initialisation of variables differently.

// In SystemVerilog, initialisation happens before
// any events and does itself not cause any events
// to happen.

// So, e.g. the following will always print 0:

logic a = 0;

initial $display("a = %b", a);

// In Verilog before SystemVerilog, the above
// had the following semantics
// (with "a" renamed to "b"):

logic b;

initial b = 0;

initial $display("b = %b", b);

// Which can print either x or 0, because the order
// of the initial processes is nondeterministic.

endmodule
