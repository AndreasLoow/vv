module display_empty1;

initial $display();

endmodule
