module always_comb_delay1;

logic a;

always_comb #1 a = 1;

endmodule
