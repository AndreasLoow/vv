module monitor2;

// Edge-case with only $time

initial $monitor("%d", $time);

endmodule
