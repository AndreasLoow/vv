module cont_var3;

// Alternative order, see cont_var2

logic a;

assign a = 1;

always @(*) a = 0;

endmodule
