module display;

initial $display("%b", $time);

endmodule
