module final1;

logic a;

// Final blocks are run after simulation has ended

final a = 0;

endmodule
