module monitor3;

// Another edge-case, with only $time

initial $monitor("%d", $time);

endmodule
