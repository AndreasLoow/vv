module monitor;

// Basic $monitor example

// (Note that the order of execution does not matter, the output is the same.)

logic a;
   
initial $monitor("a = %b at time %d", a, $time);

initial begin
 a = 1'b0;
 #10 a = 1'bz;
end

endmodule
